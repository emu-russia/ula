// Model for the classic MOSTEK 4116 16384 x 1 Bit Dynamic Ram

module MK4116 ();

endmodule // MK4116